`timescale 1ns/1ps
module float_mul_tb();
//#(parameter M = 2 ,parameter N =2,parameter P =2 )


 reg clk;
  reg reset;

  logic [0:3][31:0] a_in; // MxN matrix A
  logic [0:3][31:0] b_in; // NxP matrix B

  logic [0:3][31:0] c_out; // MxP result matrix C


fp_matrix #(.N(2), .M(2), .P(2)) uut(.clk(clk),.reset(reset), .a_in(a_in),.b_in(b_in), .c_out(c_out));

initial
begin
    clk=0;
    reset=0;
end

always #5 clk = ~clk;

initial begin

a_in = {32'b00111111100000000000000000000000, 32'b01000000000000000000000000000000,32'b01000000010000000000000000000000, 32'b01000000100000000000000000000000};
b_in = {32'b01000000101000000000000000000000, 32'b01000000110000000000000000000000,32'b01000000111000000000000000000000, 32'b01000001000000000000000000000000};

//        a_in[0][0] = 32'b01000000100000000000000000000000;//1
        
//        a_in[0][1] = 32'b01000000010000000000000000000000;//2
           
//        a_in[1][0] = 32'b01000000100000000000000000000000;//3
        
//        a_in[1][1] = 32'b01000000010000000000000000000000;//4
        
////        a_in[4] = 32'b01000000100000000000000000000000;//5.75
        
////        a_in[5] = 32'b01000000010000000000000000000000;//6.75
        

//        b_in[0][0] = 32'b01000000100000000000000000000000;//5
        
//        b_in[0][1] = 32'b01000000010000000000000000000000;//6
            
//        b_in[1][0] = 32'b01000000100000000000000000000000;//7
        
//        b_in[1][1] = 32'b01000000010000000000000000000000;//8
        
////        b_in[4] = 32'b01000000100000000000000000000000;//7.375
        
////        b_in[5] = 32'b01000000010000000000000000000000;//8.375

//        //result should be 28,21,28,21 
////01000010111111100111000000000000
////01000010111111100111000000000000

//

       
end



initial
begin

//$dumpfile("float_matrix.vcd");
//$dumpvars(0,float_mul_tb);

    #2000
    $finish;
end


endmodule